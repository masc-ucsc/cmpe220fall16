`ifndef SCMEM_H
`define SCMEM_H

`include "scmemp.vh"
`include "scmemc.vh"
`include "scmemt.vh"
`include "scmemi.vh"

`endif

