
module top_2core2dr(
   input                           clk
  ,input                           reset
);

 // net_2core2dr
 // L1, L2, DR
 //
 // In/out: L1 interface, pfengine, directory_memory requests

endmodule

